module nonresdiv(D, R_0, Q, R_n1);
  input [1:0] D;
  output [2:0] Q;
  input [3:0] R_0;
  output [4:0] R_n1;
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  assign _000_ = R_0[3] & ~(D[1]);
  assign _001_ = R_0[2] | ~(D[0]);
  assign _002_ = R_0[3] ^ D[1];
  assign _003_ = _001_ & ~(_002_);
  assign _004_ = ~(_003_ | _000_);
  assign Q[2] = ~_004_;
  assign _005_ = ~D[1];
  assign _006_ = _004_ ^ _005_;
  assign _007_ = ~(R_0[2] ^ D[0]);
  assign _008_ = _006_ & ~(_007_);
  assign _009_ = _004_ ^ D[0];
  assign _010_ = R_0[1] & ~(_009_);
  assign _011_ = ~R_0[0];
  assign _012_ = _011_ & ~(_004_);
  assign _013_ = R_0[0] & ~(_004_);
  assign _014_ = _013_ | _012_;
  assign _015_ = _009_ ^ R_0[1];
  assign _016_ = _014_ & ~(_015_);
  assign _017_ = _016_ | _010_;
  assign _018_ = _007_ ^ _006_;
  assign _019_ = _017_ & ~(_018_);
  assign _020_ = _019_ | _008_;
  assign _021_ = _002_ ^ _001_;
  assign _022_ = ~(_021_ ^ _004_);
  assign _023_ = _020_ & ~(_022_);
  assign _024_ = ~(_021_ | _004_);
  assign Q[1] = _024_ | _023_;
  assign _025_ = _022_ ^ _020_;
  assign _026_ = Q[1] & ~(_025_);
  assign _027_ = R_0[1] ^ D[0];
  assign _028_ = Q[1] ^ D[1];
  assign _029_ = _028_ & _027_;
  assign _030_ = Q[1] | D[0];
  assign _031_ = D[0] & ~(R_0[0]);
  assign _032_ = _030_ & ~(_031_);
  assign _033_ = ~(_028_ ^ _027_);
  assign _034_ = _032_ & ~(_033_);
  assign _035_ = _034_ | _029_;
  assign _036_ = _018_ ^ _017_;
  assign _037_ = _036_ ^ Q[1];
  assign _038_ = _035_ & ~(_037_);
  assign _039_ = Q[1] & ~(_036_);
  assign _040_ = _039_ | _038_;
  assign _041_ = _025_ ^ Q[1];
  assign _042_ = _040_ & ~(_041_);
  assign Q[0] = _042_ | _026_;
  assign _043_ = _033_ ^ _032_;
  assign _044_ = ~_043_;
  assign _045_ = D[1] & ~(Q[0]);
  assign _046_ = ~(_045_ & _044_);
  assign _047_ = R_0[0] ^ D[0];
  assign _048_ = Q[0] | ~(D[0]);
  assign _049_ = _047_ & ~(_048_);
  assign _050_ = _045_ ^ _044_;
  assign _051_ = _050_ & _049_;
  assign _052_ = _046_ & ~(_051_);
  assign _053_ = _037_ ^ _035_;
  assign _054_ = _053_ | _052_;
  assign _055_ = _041_ ^ _040_;
  assign R_n1[3] = _055_ ^ _054_;
  assign R_n1[0] = ~(_048_ ^ _047_);
  assign R_n1[1] = _050_ ^ _049_;
  assign R_n1[2] = _053_ ^ _052_;
  assign _056_ = _055_ | _054_;
  assign R_n1[4] = _056_ ^ Q[0];
endmodule
